`include "testbench.v"
`include "decimal_display.v"

module decimal_display_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
