`include "btn_in.v"

module btn_in_tb;
endmodule
