`include "decimal_decoder.v"

module decimal_decoder_tb;
endmodule
