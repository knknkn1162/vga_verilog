`include "hex_decoder.v"

module hex_decoder_tb;
endmodule
