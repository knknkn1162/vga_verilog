`include "testbench.v"
`include "px_clk.v"

module px_clk_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
