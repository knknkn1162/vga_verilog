`include "testbench.v"
`include "top.v"

module top_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
