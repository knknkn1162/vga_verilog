`include "testbench.v"
`include "rgb.v"

module rgb_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
