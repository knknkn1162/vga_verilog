`include "testbench.v"
`include "hsync.v"

module hsync_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
