`include "testbench.v"
`include "gen_640_480.v"

module gen_640_480_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
