`include "testbench.v"
`include "hex_display.v"

module hex_display_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
