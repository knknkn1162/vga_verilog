`include "testbench.v"
`include "vsync.v"

module vsync_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
